3.5


R1 X 0 1
C1 X 0 1u ic=1.33
R2 X 3 2
V2 3 0 dc 2V
.tran 10p 10u uic

.control
set filetype=ascii
run
plot v(X)
wrdata 3.5.dat v(X)
//set gnuplot_terminal=pdf/quit
//gnuplot ../figs/3.5 v(X) 
.endc

.end